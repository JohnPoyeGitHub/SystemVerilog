input logic [2:0] a;
input logic nxt_bit;
input logic [2:0] b;
input logic [2:0] R;
output logi