module cla_8bit (
    input  logic [7:0] A,
    input  logic [7:0] B,
    output logic [8:0] Sum
);

 
endmodule
