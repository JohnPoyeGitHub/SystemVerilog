module rca_nbit #(parameter N = 4)(
	input logic [N-1:0] a,
	input logic [N-1:0] b,
	input logic cin,
	output logic [N-1:0] sum,
	output logic co
);

//
endmodule