logic input [N]a;
logic input [N]b;