logic input [N:0]a;
logic input [N:0]b;
logic output [N+1:0]y;

