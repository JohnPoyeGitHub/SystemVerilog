logic input a;
